// Project F Library - 640x480p60 Display
// (C)2022 Will Green, open source hardware released under the MIT License
// Learn more at https://projectf.io

module HDMISigGen #(
    CORDW=16,    // signed coordinate width (bits)
    H_RES=640,   // horizontal resolution (pixels)
    V_RES=480,   // vertical resolution (lines)
    H_FP=16,     // horizontal front porch
    H_SYNC=96,   // horizontal sync
    H_BP=48,     // horizontal back porch
    V_FP=10,     // vertical front porch
    V_SYNC=2,    // vertical sync
    V_BP=33,     // vertical back porch
    H_POL=0,     // horizontal sync polarity (0:neg, 1:pos)
    V_POL=0      // vertical sync polarity (0:neg, 1:pos)
)(
    input  logic                    i_clk_pix, // pixel clock 25mhz
    input  logic                    i_rst_pix, // reset in pixel clock domain
    output logic                    o_hsync,   // horizontal sync
    output logic                    o_vsync,   // vertical sync
    output logic                    o_de,      // data enable (low in blanking interval)
    output logic                    o_frame,   // high at start of frame (include prev frame blank)
    output logic                    o_line,    // high at start of line (include prev frame blank)             
    output logic signed [CORDW-1:0] o_sx,      // horizontal screen position
    output logic signed [CORDW-1:0] o_sy       // vertical screen position
);

    // horizontal timings
    localparam signed H_STA  = 0 - H_FP - H_SYNC - H_BP;    // horizontal start
    localparam signed HS_STA = H_STA + H_FP;                // sync start
    localparam signed HS_END = HS_STA + H_SYNC;             // sync end
    localparam signed HA_STA = 0;                           // active start
    localparam signed HA_END = H_RES - 1;                   // active end

    // vertical timings
    localparam signed V_STA  = 0 - V_FP - V_SYNC - V_BP;    // vertical start
    localparam signed VS_STA = V_STA + V_FP;                // sync start
    localparam signed VS_END = VS_STA + V_SYNC;             // sync end
    localparam signed VA_STA = 0;                           // active start
    localparam signed VA_END = V_RES - 1;                   // active end

    logic signed [CORDW-1:0] x, y;  // screen position

    // generate horizontal and vertical sync with correct polarity
    always_ff @(posedge i_clk_pix) begin
        o_hsync <= H_POL ? (x > HS_STA && x <= HS_END) : ~(x > HS_STA && x <= HS_END);
        o_vsync <= V_POL ? (y > VS_STA && y <= VS_END) : ~(y > VS_STA && y <= VS_END);
        if (i_rst_pix) begin
            o_hsync <= H_POL ? 0 : 1;
            o_vsync <= V_POL ? 0 : 1;
        end
    end

    // control signals
    always_ff @(posedge i_clk_pix) begin
        o_de    <= (y >= VA_STA && x >= HA_STA);
        o_frame <= (y == V_STA  && x == H_STA);
        o_line  <= (x == H_STA);
        if (i_rst_pix) begin
            o_de <= 0;
            o_frame <= 0;
            o_line <= 0;
        end
    end

    // calculate horizontal and vertical screen position
    always_ff @(posedge i_clk_pix) begin
        if (x == HA_END) begin  // last pixel on o_line?
            x <= H_STA;
            y <= (y == VA_END) ? V_STA : y + 1;  // last o_line on screen?
        end else begin
            x <= x + 1;
        end
        if (i_rst_pix) begin
            x <= H_STA;
            y <= V_STA;
        end
    end

    // delay screen position to match sync and control signals
    always_ff @ (posedge i_clk_pix) begin
        o_sx <= x;
        o_sy <= y;
        if (i_rst_pix) begin
            o_sx <= H_STA;
            o_sy <= V_STA;
        end
    end
endmodule
